module easy_verilog_example(

    );
	
	reg x = 1'b0; // 1bit variable with the value 0
	reg y = 1'b1; // 1bit variable with the value 1	
	reg z;        // used to store the result of operations between x and y

    // A procedure example
    always @(*) begin
        $display("x=%b, y=%b, z=%b", x,y,z);
	end
	
	// Another procedure example
	initial begin
        #2;         // wait 2 time units
        z = x ^ y;  // bit-wise XOR between the 1 bit variables x and y    
	    #10;        // wait 10 time units
        y = 0;      // change the value of y
        z = x | y;  // bit-wise OR between the 1 bit variables x and y   
        #10;        // wait 10 time units
        z = z & 1;  // bit-wise AND between the 1 bit variable z and 1
        #10;        // wait 10 time units
	end

endmodule{"threads":[{"position":415,"start":0,"end":414,"connection":"closed"},{"position":415,"start":415,"end":828,"connection":"open"}],"url":"https://att-c.udemycdn.com/2021-08-26_13-58-14-eef4e0f315fd039da49d90ad6a823394/original.v?response-content-disposition=attachment%3B+filename%3Deasy_verilog_example.v&Expires=1632531454&Signature=aBuxkdRrSVGNDetOEfa~vVhYA4Bj8bBaRY7Q69YVEEmDrZ3krQw~FcMfSH1sdUfZrQ5MSd279XmQdOYTmemWChHSshMxOwFHBPgG19Gcn7SfOqReWDhyLEwdm2UG6B4OqRAsnP21cZPNqMYqEVpfkLT0H2OK30BGEa2o5KvYNji1lh~vXHuZedMJ-9CTWimmxY-a~EOZSPeZY0OQFHa1Gx9yjbrGa1u~aMxqpT8er0FCaqJy9IbLcnnfvzLSG6GELNjuXeeaIsMrQoUz5aMfDLzu0f0a1VQyVshmzTbsut1pCYEnL2PtJ~3f48cSoncmy-cgt~QlLS~eL~vab4kF0w__&Key-Pair-Id=APKAITJV77WS5ZT7262A","method":"GET","port":443,"downloadSize":828,"headers":{"content-type":"binary/octet-stream","content-length":"828","connection":"close","date":"Fri, 24 Sep 2021 20:28:00 GMT","last-modified":"Thu, 26 Aug 2021 13:58:17 GMT","etag":"\"381a3ae89bfb960e71d90cbd03dfd740\"","x-amz-server-side-encryption":"AES256","x-amz-meta-qqfilename":"easy_verilog_example.v","x-amz-version-id":"LWxDKsLcaEip2uimEdKrMyPLBvPpmttK","content-disposition":"attachment; filename=easy_verilog_example.v","accept-ranges":"bytes","server":"AmazonS3","x-edge-origin-shield-skipped":"0, 0","x-cache":"Miss from cloudfront","via":"1.1 e0efba8a72628bfc3dc6d4d637b28302.cloudfront.net (CloudFront)","x-amz-cf-pop":"FRA2-C1","x-amz-cf-id":"llTLHDkrUA4PsWZ9Gjx-136AsrcgV_t-MrMBV1RU3NQYvXcK7KurbQ=="}}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      