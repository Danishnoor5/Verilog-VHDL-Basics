module prio_enc2_4to2
  (input [3:0] d,
   output reg [1:0] q,
   output reg v
  );
  
    always @(*) begin
        case (1) // checks if a signal is set
            d[3]:  begin q = 2'd3; v = 1; end
            d[2]:  begin q = 2'd2; v = 1; end
            d[1]:  begin q = 2'd1; v = 1; end
            d[0]:  begin q = 2'd0; v = 1; end
            default: begin q = 2'd0; v = 0; end
        endcase
    end
  
endmodule


`timescale 1us/1ns
module tb_prio_enc2_4to2();
	
    reg [3:0] d;   // DUT variables
    wire v;
    wire [1:0] q;
    integer i;     // testbench variable

    // Instantiate the DUT 
    prio_enc2_4to2 PRENC(
      .d(d),
      .q(q),
      .v(v)
    );
  
    // Create stimulus
    initial begin
        $monitor($time, " d = %b, q = %d, v = %d", d, q, v);
        #1; d = 0; 
        for (i = 0; i<4; i=i+1) begin
           #1; d = (1 << i);
        end
        #1; d = 4'b1111;
        #1; d = 4'b1001;
        #1; d = 4'b0101;
		#1; d = 4'b0000;
		#1; $stop;
    end
  
endmodule
{"threads":[{"position":533,"start":0,"end":532,"connection":"closed"},{"position":533,"start":533,"end":1063,"connection":"open"}],"url":"https://att-c.udemycdn.com/2021-08-30_12-53-16-58bb20c70ded4f93902b7dfbc59920f2/original.v?response-content-disposition=attachment%3B+filename%3Dprio_enc2_4to2.v&Expires=1632531454&Signature=YtDlXC9UPYLF8BdoKMmtEJxJr2-WrgjAVpx8vT4TRn0OZg7qRjedVBk5IZDJXQq9hdkSbkLt9kBNllc4tBDziXvXWZwxjHgVOcBjmz~ncVRJ4pJOFCtpXYbnTIMe84tyUnHg2t7a00SAlSN4FhYggcZ9MaUJk0-qe7R2yXFeb2LHrBGgsZh2J2QZ9g8hxTOFHKy~pcLK-iPPdSouIo2TN8O59StjvY5540fCVXE3dJNkaNkOqgjb7FQl1JSQTyCe97iSiIgqpvE3Z~kpMeiqfoS54nTtpfmcL7wMaPGCh5SVWdN5DQCUDMsN00z~LPIfl6asUf4xX-RcjexoAC3zMw__&Key-Pair-Id=APKAITJV77WS5ZT7262A","method":"GET","port":443,"downloadSize":1063,"headers":{"content-type":"binary/octet-stream","content-length":"1063","connection":"close","date":"Fri, 24 Sep 2021 20:30:32 GMT","last-modified":"Mon, 30 Aug 2021 12:53:17 GMT","etag":"\"4767c5b38484552241f74dc31ad2b820\"","x-amz-server-side-encryption":"AES256","x-amz-meta-qqfilename":"prio_enc2_4to2.v","x-amz-version-id":"xtcRaVpKA3jiX.I2s5xJtANE8st6luNk","content-disposition":"attachment; filename=prio_enc2_4to2.v","accept-ranges":"bytes","server":"AmazonS3","x-edge-origin-shield-skipped":"0, 0","x-cache":"Miss from cloudfront","via":"1.1 69f13f852a135432abb1b7bfc5a8b421.cloudfront.net (CloudFront)","x-amz-cf-pop":"FRA2-C1","x-amz-cf-id":"cdZHojJG0hptn6EYuZp6Lwd9CQUH1WKF9c8j1zsxF83hmN1QKcUiBQ=="}}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     